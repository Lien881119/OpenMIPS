`include "define.v"
`include "openmips_min_sopc.v"
`timescale 1ns/1ps

module openmips_min_sopc_tb();

    initial
    begin            
        $dumpfile("wave.vcd");        
        $dumpvars(0, openmips_min_sopc_tb);
    end
    reg CLOCK_50;
    reg rst;

    initial begin
        CLOCK_50 = 1'b0;
        forever #10 CLOCK_50 = ~CLOCK_50;
    end

    initial begin
        rst = `RstEnable;
        #195 rst = `RstDisable;
        #1000 $stop;
    end

    //initialize sopc
    openmips_min_sopc openmips_min_sopc0(.clk(CLOCK_50), .rst(rst));

endmodule