`include "define.v"

module id_ex (
    input wire clk,
    input wire rst,
);
    
endmodule